.title KiCad schematic
V1 /IN 0 AC 1
R1 /OUT /IN {RLPF}
C1 /OUT 0 {CLPF}
.end
